mynetlist
R1 6 1 100
R2 1 0 100
R3 1 2 100 
R4 2 3 100
R5 3 0 100
R6 2 5 100
R7 5 0 100
.control
op
print v(1) v(2) v(3) v(4) v(5) v(6) 
.endc
.end
