mynetlist
Vt4 4 0 DC 1
Vg1 1 0 DC 0
Vg2 2 0 DC 0
R0 1 2 92
R1 1 3 17
R2 1 4 88
R3 2 3 56
R4 3 4 84
R5 4 0 81
.control
    op
    print v(1) v(2) v(3) v(4) 
print i(Vt4)
    .endc
    .end
    